`define DSIZE 8
//`define ASIZE $clog2(`DSIZE)
`define ASIZE 3
`define no_of_trxn 100
