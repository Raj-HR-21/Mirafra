`include "defines.sv"

package alu_pkg;

`include "alu_transaction.sv"
`include "alu_generator.sv"
`include "alu_driver.sv"
`include "alu_monitor.sv"
`include "alu_ref_model.sv"
`include "alu_scb.sv"
`include "alu_env.sv"
`include "alu_test.sv"

endpackage
