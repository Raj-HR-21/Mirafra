
package alu_pkg;
`include "uvm_pkg.sv"
`include "uvm_macros.svh"
	import uvm_pkg::*;
	`include "seq_item.sv"
	`include "sequence.sv"
	`include "sequencer.sv"
	`include "driver.sv"
	`include "monitor.sv"
	`include "agent.sv"
	`include "scoreboard.sv"
	`include "subscriber.sv"
	`include "env.sv"
	`include "test.sv"


endpackage
